`timescale 1ns / 1ns

module wave_generator(
    input wire clk,
    input wire [15:0] freq,
    output reg signed [9:0] wave_out
);
    reg [5:0] i;
    reg signed [7:0] amplitude [0:63];
    reg [15:0] counter = 0;

    initial begin
        amplitude[0] = 0;
        amplitude[1] = 7;
        amplitude[2] = 13;
        amplitude[3] = 19;
        amplitude[4] = 25;
        amplitude[5] = 30;
        amplitude[6] = 35;
        amplitude[7] = 40;
        amplitude[8] = 45;
        amplitude[9] = 49;
        amplitude[10] = 52;
        amplitude[11] = 55;
        amplitude[12] = 58;
        amplitude[13] = 60;
        amplitude[14] = 62;
        amplitude[15] = 63;
        amplitude[16] = 63;
        amplitude[17] = 63;
        amplitude[18] = 62;
        amplitude[19] = 60;
        amplitude[20] = 58;
        amplitude[21] = 55;
        amplitude[22] = 52;
        amplitude[23] = 49;
        amplitude[24] = 45;
        amplitude[25] = 40;
        amplitude[26] = 35;
        amplitude[27] = 30;
        amplitude[28] = 25;
        amplitude[29] = 19;
        amplitude[30] = 13;
        amplitude[31] = 7;
        amplitude[32] = 0;
        amplitude[33] = -7;
        amplitude[34] = -13;
        amplitude[35] = -19;
        amplitude[36] = -25;
        amplitude[37] = -30;
        amplitude[38] = -35;
        amplitude[39] = -40;
        amplitude[40] = -45;
        amplitude[41] = -49;
        amplitude[42] = -52;
        amplitude[43] = -55;
        amplitude[44] = -58;
        amplitude[45] = -60;
        amplitude[46] = -62;
        amplitude[47] = -63;
        amplitude[48] = -63;
        amplitude[49] = -63;
        amplitude[50] = -62;
        amplitude[51] = -60;
        amplitude[52] = -58;
        amplitude[53] = -55;
        amplitude[54] = -52;
        amplitude[55] = -49;
        amplitude[56] = -45;
        amplitude[57] = -40;
        amplitude[58] = -35;
        amplitude[59] = -30;
        amplitude[60] = -25;
        amplitude[61] = -19;
        amplitude[62] = -13;
        amplitude[63] = -7;
    end

    always @ (posedge clk) begin
      if (freq == 0) wave_out <= 0;
      else
      if (counter == freq) begin
        counter <= 0;
        wave_out <= $signed(amplitude[i]);
        i <= i + 1;
        if (i == 63) i <= 0; else i <= i + 1;
      end else counter <= counter + 1;
    end
endmodule

module audio_output(
  input wire clk,
  output reg out
);
    wire signed [9:0] ch[0:4];
    wire signed [11:0] wave_sum;
    wire [11:0] positive_wave_sum;
    wire [15:0] freq_count [0:4];
    reg [9:0] PWM;
    reg [31:0] music_data [0:79];
    reg [31:0] music_data2 [0:79];
    reg [31:0] music_data3 [0:180];
    reg [31:0] play_counter;
    reg [15:0] note_counter = 0;
    reg [15:0] note_counter1 = 0;
    reg [31:0] note_data[0:1];
    reg [31:0] note_data2;
    wave_generator ch0(clk, freq_count[0], ch[0]);
    wave_generator ch1(clk, freq_count[1], ch[1]);
    wave_generator ch2(clk, freq_count[2], ch[2]);
    assign freq_count[0] = note_data[0][31:16];
    assign freq_count[1] = note_data[1][31:16];
    assign freq_count[2] = note_data2[31:16];
    assign wave_sum = ch[2] + ch[1] + ch[0];
    assign positive_wave_sum = wave_sum * 2 + 512;
    initial begin
    music_data[0] = 32'h0000010a;
    music_data[1] = 32'h1284010a;
    music_data[2] = 32'h1754010a;
    music_data[3] = 32'h18b7010a;
    music_data[4] = 32'h0ddf010a;
    music_data[5] = 32'h0d17010a;
    music_data[6] = 32'h14c80085;
    music_data[7] = 32'h0c5b0085;
    music_data[8] = 32'h14c80085;
    music_data[9] = 32'h00000085;
    music_data[10] = 32'h0c5b0085;
    music_data[11] = 32'h00000085;
    music_data[12] = 32'h0c5b0215;
    music_data[13] = 32'h0000010a;
    music_data[14] = 32'h0f91026e;
    music_data[15] = 32'h000000b1;
    music_data[16] = 32'h107f026e;
    music_data[17] = 32'h000000b1;
    music_data[18] = 32'h0f91026e;
    music_data[19] = 32'h00000137;
    music_data[20] = 32'h00000085;
    music_data[21] = 32'h00000085;
    music_data[22] = 32'h00000085;
    music_data[23] = 32'h00000085;
    music_data[24] = 32'h00000085;
    music_data[25] = 32'h0f91026e;
    music_data[26] = 32'h000000b1;
    music_data[27] = 32'h107f0215;
    music_data[28] = 32'h08bd010a;
    music_data[29] = 32'h0f91026e;
    music_data[30] = 32'h0000034c;
    music_data[31] = 32'h00000085;
    music_data[32] = 32'h117a026e;
    music_data[33] = 32'h000000b1;
    music_data[34] = 32'h0b02026e;
    music_data[35] = 32'h000000b1;
    music_data[36] = 32'h117a026e;
    music_data[37] = 32'h00000137;
    music_data[38] = 32'h00000085;
    music_data[39] = 32'h00000085;
    music_data[40] = 32'h00000085;
    music_data[41] = 32'h00000085;
    music_data[42] = 32'h00000085;
    music_data[43] = 32'h0a64026e;
    music_data[44] = 32'h000000b1;
    music_data[45] = 32'h0f910215;
    music_data[46] = 32'h0ddf010a;
    music_data[47] = 32'h0f91026e;
    music_data[48] = 32'h0000034c;
    music_data[49] = 32'h00000085;
    music_data[50] = 32'h0942026e;
    music_data[51] = 32'h000000b1;
    music_data[52] = 32'h07c8026e;
    music_data[53] = 32'h000000b1;
    music_data[54] = 32'h07c8026e;
    music_data[55] = 32'h000000b1;
    music_data[56] = 32'h0000010a;
    music_data[57] = 32'h00000085;
    music_data[58] = 32'h0000010a;
    music_data[59] = 32'h00000085;
    music_data[60] = 32'h08bd026e;
    music_data[61] = 32'h000000b1;
    music_data[62] = 32'h08bd026e;
    music_data[63] = 32'h000000b1;
    music_data[64] = 32'h0baa026e;
    music_data[65] = 32'h000000b1;
    music_data[66] = 32'h0000010a;
    music_data[67] = 32'h00000085;
    music_data[68] = 32'h0000010a;
    music_data[69] = 32'h00000085;
    music_data[70] = 32'h0942026e;
    music_data[71] = 32'h000000b1;
    music_data[72] = 32'h117a010a;
    music_data[73] = 32'h0c5b010a;
    music_data[74] = 32'h0c5b010a;
    music_data[75] = 32'h09420085;
    music_data[76] = 32'h0c5b0085;
    music_data[77] = 32'h0942018f;
    music_data[78] = 32'h117a0085;
    music_data[79] = 32'h1284031f;
    music_data2[0] = 32'h14c8010a;
    music_data2[1] = 32'h1605010a;
    music_data2[2] = 32'h107f010a;
    music_data2[3] = 32'h0f91010a;
    music_data2[4] = 32'h1754010a;
    music_data2[5] = 32'h1605010a;
    music_data2[6] = 32'h0c5b0085;
    music_data2[7] = 32'h14c80085;
    music_data2[8] = 32'h0c5b0085;
    music_data2[9] = 32'h00000085;
    music_data2[10] = 32'h12840085;
    music_data2[11] = 32'h00000085;
    music_data2[12] = 32'h117a0215;
    music_data2[13] = 32'h0f91010a;
    music_data2[14] = 32'h0942026e;
    music_data2[15] = 32'h000000b1;
    music_data2[16] = 32'h09cf026e;
    music_data2[17] = 32'h000000b1;
    music_data2[18] = 32'h0942026e;
    music_data2[19] = 32'h00000137;
    music_data2[20] = 32'h0f910085;
    music_data2[21] = 32'h0ddf0085;
    music_data2[22] = 32'h0c5b0085;
    music_data2[23] = 32'h0baa0085;
    music_data2[24] = 32'h0a640085;
    music_data2[25] = 32'h0942026e;
    music_data2[26] = 32'h000000b1;
    music_data2[27] = 32'h09cf0215;
    music_data2[28] = 32'h0ddf010a;
    music_data2[29] = 32'h0942026e;
    music_data2[30] = 32'h0000034c;
    music_data2[31] = 32'h0f910085;
    music_data2[32] = 32'h0a64026e;
    music_data2[33] = 32'h000000b1;
    music_data2[34] = 32'h1284026e;
    music_data2[35] = 32'h000000b1;
    music_data2[36] = 32'h0a64026e;
    music_data2[37] = 32'h00000137;
    music_data2[38] = 32'h0f910085;
    music_data2[39] = 32'h0ddf0085;
    music_data2[40] = 32'h0c5b0085;
    music_data2[41] = 32'h0baa0085;
    music_data2[42] = 32'h0b020085;
    music_data2[43] = 32'h117a026e;
    music_data2[44] = 32'h000000b1;
    music_data2[45] = 32'h18b70215;
    music_data2[46] = 32'h08bd010a;
    music_data2[47] = 32'h0942026e;
    music_data2[48] = 32'h0000034c;
    music_data2[49] = 32'h0f910085;
    music_data2[50] = 32'h07c8026e;
    music_data2[51] = 32'h000000b1;
    music_data2[52] = 32'h0a64026e;
    music_data2[53] = 32'h000000b1;
    music_data2[54] = 32'h0b02026e;
    music_data2[55] = 32'h000000b1;
    music_data2[56] = 32'h07c8010a;
    music_data2[57] = 32'h06ef0085;
    music_data2[58] = 32'h0000010a;
    music_data2[59] = 32'h07c80085;
    music_data2[60] = 32'h0a64026e;
    music_data2[61] = 32'h000000b1;
    music_data2[62] = 32'h0b02026e;
    music_data2[63] = 32'h000000b1;
    music_data2[64] = 32'h08bd026e;
    music_data2[65] = 32'h000000b1;
    music_data2[66] = 32'h08bd010a;
    music_data2[67] = 32'h07c80085;
    music_data2[68] = 32'h0000010a;
    music_data2[69] = 32'h08bd0085;
    music_data2[70] = 32'h1754026e;
    music_data2[71] = 32'h000000b1;
    music_data2[72] = 32'h0ddf010a;
    music_data2[73] = 32'h0f91010a;
    music_data2[74] = 32'h08bd010a;
    music_data2[75] = 32'h0c5b0085;
    music_data2[76] = 32'h09420085;
    music_data2[77] = 32'h0c5b018f;
    music_data2[78] = 32'h0c5b0085;
    music_data2[79] = 32'h0baa031f;
    music_data3[0] = 32'h00000855;
    music_data3[1] = 32'h1f230085;
    music_data3[2] = 32'h00000085;
    music_data3[3] = 32'h1f23031f;
    music_data3[4] = 32'h2ea80085;
    music_data3[5] = 32'h00000085;
    music_data3[6] = 32'h1f230085;
    music_data3[7] = 32'h00000085;
    music_data3[8] = 32'h17540085;
    music_data3[9] = 32'h00000085;
    music_data3[10] = 32'h316e0085;
    music_data3[11] = 32'h00000085;
    music_data3[12] = 32'h1f230085;
    music_data3[13] = 32'h00000085;
    music_data3[14] = 32'h18b70085;
    music_data3[15] = 32'h00000085;
    music_data3[16] = 32'h2ea80085;
    music_data3[17] = 32'h00000085;
    music_data3[18] = 32'h1f230085;
    music_data3[19] = 32'h00000085;
    music_data3[20] = 32'h17540085;
    music_data3[21] = 32'h00000085;
    music_data3[22] = 32'h25080085;
    music_data3[23] = 32'h00000085;
    music_data3[24] = 32'h1f230085;
    music_data3[25] = 32'h00000085;
    music_data3[26] = 32'h17540085;
    music_data3[27] = 32'h00000085;
    music_data3[28] = 32'h2ea80085;
    music_data3[29] = 32'h00000085;
    music_data3[30] = 32'h1f230085;
    music_data3[31] = 32'h00000085;
    music_data3[32] = 32'h17540085;
    music_data3[33] = 32'h00000085;
    music_data3[34] = 32'h316e0085;
    music_data3[35] = 32'h00000085;
    music_data3[36] = 32'h1f230085;
    music_data3[37] = 32'h00000085;
    music_data3[38] = 32'h18b70085;
    music_data3[39] = 32'h00000085;
    music_data3[40] = 32'h2ea80085;
    music_data3[41] = 32'h00000085;
    music_data3[42] = 32'h1f230085;
    music_data3[43] = 32'h00000085;
    music_data3[44] = 32'h17540085;
    music_data3[45] = 32'h00000085;
    music_data3[46] = 32'h25080085;
    music_data3[47] = 32'h00000085;
    music_data3[48] = 32'h1f230085;
    music_data3[49] = 32'h00000085;
    music_data3[50] = 32'h17540085;
    music_data3[51] = 32'h00000085;
    music_data3[52] = 32'h29910085;
    music_data3[53] = 32'h00000085;
    music_data3[54] = 32'h1f230085;
    music_data3[55] = 32'h00000085;
    music_data3[56] = 32'h18b70085;
    music_data3[57] = 32'h00000085;
    music_data3[58] = 32'h2c0a0085;
    music_data3[59] = 32'h00000085;
    music_data3[60] = 32'h20fe0085;
    music_data3[61] = 32'h00000085;
    music_data3[62] = 32'h1a2f0085;
    music_data3[63] = 32'h00000085;
    music_data3[64] = 32'h29910085;
    music_data3[65] = 32'h00000085;
    music_data3[66] = 32'h1f230085;
    music_data3[67] = 32'h00000085;
    music_data3[68] = 32'h18b70085;
    music_data3[69] = 32'h00000085;
    music_data3[70] = 32'h316e0085;
    music_data3[71] = 32'h00000085;
    music_data3[72] = 32'h1f230085;
    music_data3[73] = 32'h00000085;
    music_data3[74] = 32'h18b70085;
    music_data3[75] = 32'h00000085;
    music_data3[76] = 32'h29910085;
    music_data3[77] = 32'h00000085;
    music_data3[78] = 32'h1f230085;
    music_data3[79] = 32'h00000085;
    music_data3[80] = 32'h18b70085;
    music_data3[81] = 32'h00000085;
    music_data3[82] = 32'h316e0085;
    music_data3[83] = 32'h00000085;
    music_data3[84] = 32'h1f230085;
    music_data3[85] = 32'h00000085;
    music_data3[86] = 32'h18b70085;
    music_data3[87] = 32'h00000085;
    music_data3[88] = 32'h2ea80085;
    music_data3[89] = 32'h00000085;
    music_data3[90] = 32'h1f230085;
    music_data3[91] = 32'h00000085;
    music_data3[92] = 32'h17540085;
    music_data3[93] = 32'h00000085;
    music_data3[94] = 32'h3e470085;
    music_data3[95] = 32'h00000085;
    music_data3[96] = 32'h1f230085;
    music_data3[97] = 32'h00000085;
    music_data3[98] = 32'h17540085;
    music_data3[99] = 32'h00000085;
    music_data3[100] = 32'h2ea80085;
    music_data3[101] = 32'h00000085;
    music_data3[102] = 32'h1f230085;
    music_data3[103] = 32'h00000085;
    music_data3[104] = 32'h12840085;
    music_data3[105] = 32'h00000085;
    music_data3[106] = 32'h316e0085;
    music_data3[107] = 32'h00000085;
    music_data3[108] = 32'h1f230085;
    music_data3[109] = 32'h00000085;
    music_data3[110] = 32'h14c80085;
    music_data3[111] = 32'h00000085;
    music_data3[112] = 32'h345f0085;
    music_data3[113] = 32'h00000085;
    music_data3[114] = 32'h1f230085;
    music_data3[115] = 32'h00000085;
    music_data3[116] = 32'h16050085;
    music_data3[117] = 32'h00000085;
    music_data3[118] = 32'h2c0a0085;
    music_data3[119] = 32'h00000085;
    music_data3[120] = 32'h1f230085;
    music_data3[121] = 32'h00000085;
    music_data3[122] = 32'h12840085;
    music_data3[123] = 32'h00000085;
    music_data3[124] = 32'h29910085;
    music_data3[125] = 32'h00000085;
    music_data3[126] = 32'h1bbe0085;
    music_data3[127] = 32'h00000085;
    music_data3[128] = 32'h117a0085;
    music_data3[129] = 32'h00000085;
    music_data3[130] = 32'h2c0a0085;
    music_data3[131] = 32'h00000085;
    music_data3[132] = 32'h1bbe0085;
    music_data3[133] = 32'h00000085;
    music_data3[134] = 32'h117a0085;
    music_data3[135] = 32'h00000085;
    music_data3[136] = 32'h2ea80085;
    music_data3[137] = 32'h00000085;
    music_data3[138] = 32'h1bbe0085;
    music_data3[139] = 32'h00000085;
    music_data3[140] = 32'h117a0085;
    music_data3[141] = 32'h00000085;
    music_data3[142] = 32'h316e0085;
    music_data3[143] = 32'h00000085;
    music_data3[144] = 32'h1f230085;
    music_data3[145] = 32'h00000085;
    music_data3[146] = 32'h117a0085;
    music_data3[147] = 32'h00000085;
    music_data3[148] = 32'h2ea80085;
    music_data3[149] = 32'h00000085;
    music_data3[150] = 32'h1f230085;
    music_data3[151] = 32'h00000085;
    music_data3[152] = 32'h12840085;
    music_data3[153] = 32'h00000085;
    music_data3[154] = 32'h3e470085;
    music_data3[155] = 32'h00000085;
    music_data3[156] = 32'h1f230085;
    music_data3[157] = 32'h00000085;
    music_data3[158] = 32'h1f230085;
    music_data3[159] = 32'h00000085;
    music_data3[160] = 32'h22f40085;
    music_data3[161] = 32'h22f40085;
    music_data3[162] = 32'h22f4018f;
    music_data3[163] = 32'h316e0085;
    music_data3[164] = 32'h2ea8031f;

    end
        parameter NOTES = 80;
        parameter BASS = 9'd165;
        parameter PLAY_DELAY = 100_000 - 1;
    always @ (posedge clk) begin
         if (play_counter == PLAY_DELAY) begin
           play_counter <= 0; 
           if (note_data2[15:0] == 0) begin
                   if (note_counter1 == BASS | note_counter1 == 0) begin note_counter1 <= 1; 
                      note_data2 <= music_data3[0]; 
                      note_counter <= 1;  note_data[0] <= music_data[0];  note_data[1] <= music_data2[0];
                      end
                   else begin note_counter1 <= note_counter1 + 1;
                      note_data2 <= music_data3[note_counter1]; 
                      end
                   end else note_data2[15:0] <= note_data2[15:0] - 1; 
           if (note_data[0][15:0] == 0) begin
               if (note_counter == 0) begin note_counter <= 1;  note_data[0] <= music_data[0];  note_data[1] <= music_data2[0];end
               else if (note_counter < NOTES) begin note_counter <= note_counter + 1; note_data[0] <= music_data[note_counter];  note_data[1] <= music_data2[note_counter]; end
           end else note_data[0][15:0] <= note_data[0][15:0] - 1;
           
         end else play_counter <= play_counter + 1; 
        if (PWM < $unsigned(positive_wave_sum)) out <= 1;
        else out <= 0;
        PWM <= PWM + 1;
    end
endmodule
/*
    set_property PACKAGE_PIN N1 [get_ports {output}]                
    set_property IOSTANDARD LVCMOS33 [get_ports {output}]
*/